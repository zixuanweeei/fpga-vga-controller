library verilog;
use verilog.vl_types.all;
entity vga_top_vga_top_sch_tb is
end vga_top_vga_top_sch_tb;
